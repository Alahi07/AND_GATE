// Code your design here
module andgate(
  input a,b,
  output y);
  assign y= a & b;
endmodule
